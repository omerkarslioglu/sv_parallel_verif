import type_pkg::*;

module task_lvl;
  
endmodule